module m_top();
  initial #200 $display("Hello, World!");
  initial begin
    #100 $display("in Verilog HDL");
    #150 $display("When am I displayed?");
  end
endmodule
