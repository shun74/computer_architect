module m_top();
  initial #200 $display("Hello, World!");
  initial #100 $display("in Verilog HDL");
endmodule
