module m_top();
  initial $display("Hello, World!");
endmodule
