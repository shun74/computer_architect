module m_top();
  initial begin
    $display("Hello, World!");
    $display("in Verilog HDL");
  end
endmodule
